pll_x14d5_inst : pll_x14d5 PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
